* NGSPICE file created from ina_top.ext - technology: sky130A

.subckt ina_top VO2 VI_2A VI_2B VI_1B VI_1A IREF VCM VO1 AVDD AVSS
X0 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 a_13371_n9266# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X4 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X5 VB2 VB2 a_22576_n12663# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X6 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X7 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X8 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X9 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X10 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X11 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X12 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X13 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X14 AVDD VB1 a_15629_n15210# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X15 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X16 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X17 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X18 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X19 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X20 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X21 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X22 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X23 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X24 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X25 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X27 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X28 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X29 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X30 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X31 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X32 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X33 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X34 AVDD VB1 a_14597_n10774# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X35 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X36 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X37 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X38 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X39 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X40 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X41 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X42 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X43 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X44 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X45 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X46 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X47 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X48 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X49 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X50 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X51 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X52 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X53 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X54 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X55 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X56 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X57 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X58 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X59 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X60 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X61 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X62 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X63 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X64 AVDD VB1 a_13887_n17331# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X65 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X66 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X67 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X68 VB4 VB4 a_22662_n9018# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X69 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X70 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X71 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X72 a_16339_n14323# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X73 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X74 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X75 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X76 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X77 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X78 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X79 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X80 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X81 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X82 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X83 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X84 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X85 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X86 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X87 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X88 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X89 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X90 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X91 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X92 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X93 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X94 VO2 VB3 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X95 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X96 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X97 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X98 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X99 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X100 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X101 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X102 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X103 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X104 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X105 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X106 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X107 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X108 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X109 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X110 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X111 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X112 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X113 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X114 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X115 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X116 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X117 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X118 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X119 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X120 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X121 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X122 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X123 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X124 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X125 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X126 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X127 a_16855_n16714# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X128 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X129 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X130 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X131 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X132 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X133 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X134 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X135 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X136 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X137 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X138 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X139 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X140 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X141 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X142 a_13887_n10774# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X143 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X144 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X145 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X146 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X147 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X148 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X149 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X150 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X151 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X152 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X153 AVSS IREF a_21723_n12663# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X154 VO1 VB3 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X155 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X156 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X157 AVDD VB1 a_14597_n13704# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X158 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X159 dda_0.VCMFB VCM dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X160 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X161 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X162 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X163 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X164 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X165 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X166 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X167 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X168 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X169 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X170 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X171 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X172 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X173 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X174 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X175 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X176 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X177 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X178 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X179 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X180 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X181 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X182 a_22662_n7484# VB4 a_22404_n7484# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X183 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X184 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X185 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X186 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X187 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X188 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X189 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X190 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X191 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X192 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X193 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X194 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X195 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X196 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X197 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X198 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X199 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X200 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X201 AVDD VB1 a_16855_n9266# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X202 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X203 AVSS IREF a_23429_n12663# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X204 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X205 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X206 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X207 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X208 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X209 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X210 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X211 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X212 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X213 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X214 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X215 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X216 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X217 a_13371_n12143# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X218 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X219 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X220 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X221 VB1 VB1 a_16339_n11522# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X222 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X223 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X224 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X225 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X226 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X227 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X228 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X229 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X230 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X231 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X232 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X233 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X234 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X235 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X236 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X237 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X238 AVDD VB1 a_14597_n15827# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X239 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X240 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X241 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X242 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X243 a_15113_n14323# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X244 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X245 VO2 VB3 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X246 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X247 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X248 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X249 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X250 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X251 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X252 AVDD VB1 a_15629_n16714# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X253 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X254 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X255 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X256 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X257 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X258 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X259 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X260 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X261 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X262 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X263 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X264 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X265 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X266 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X267 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X268 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X269 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X270 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X271 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X272 a_13887_n13704# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X273 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X274 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X275 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X276 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X277 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X278 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X279 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X280 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X281 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X282 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X283 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X284 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X285 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X286 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X287 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X288 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X289 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X290 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X291 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X292 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X293 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X294 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X295 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X296 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X297 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X298 dda_0.VIT_N1 VO1 dda_0.VD1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X299 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X300 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X301 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X302 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X303 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X304 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X305 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X306 VO1 VB3 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X307 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X308 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X309 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X310 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X311 dda_0.VCMFB VCM dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X312 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X313 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X314 a_16855_n13237# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X315 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X316 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X317 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X318 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X319 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X320 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X321 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X322 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X323 a_16339_n12143# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X324 a_22404_n7484# VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X325 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X326 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X327 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X328 a_22662_n7948# VB4 a_22404_n7948# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X329 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X330 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X331 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X332 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X333 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X334 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X335 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X336 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X337 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X338 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X339 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X340 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X341 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X342 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X343 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X344 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X345 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X346 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X347 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X348 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X349 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X350 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X351 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X352 IREF IREF a_22576_n13135# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X353 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X354 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X355 a_15629_n15210# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X356 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X357 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X358 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X359 dda_0.VIT_N2 VO2 dda_0.VD2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X360 a_15113_n9266# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X361 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X362 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X363 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X364 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X365 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X366 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X367 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X368 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X369 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X370 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X371 dda_0.VCMFB VCM dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X372 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X373 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X374 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X375 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X376 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X377 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X378 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X379 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X380 a_13887_n15827# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X381 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X382 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X383 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X384 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X385 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X386 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X387 VB3 VB1 a_15113_n10774# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X388 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X389 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X390 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X391 AVDD VB1 a_13887_n14323# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X392 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X393 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X394 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X395 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X396 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X397 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X398 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X399 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X400 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X401 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X402 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X403 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X404 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X405 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X406 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X407 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X408 AVSS IREF a_20017_n12663# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X409 dda_0.VIT_N2 VO2 dda_0.VD2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X410 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X411 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X412 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X413 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X414 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X415 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X416 dda_0.VIT_N1 VO1 dda_0.VD1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X417 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X418 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X419 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X420 VB3 VB1 a_15113_n7762# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X421 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X422 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X423 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X424 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X425 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X426 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X427 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X428 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X429 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X430 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X431 dda_0.VIT_N1 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X432 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X433 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X434 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X435 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X436 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X437 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X438 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X439 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X440 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X441 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X442 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X443 AVDD VB1 a_14597_n10153# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X444 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X445 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X446 AVDD VB1 a_15629_n13237# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X447 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X448 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X449 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X450 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X451 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X452 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X453 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X454 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X455 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X456 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X457 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X458 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X459 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X460 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X461 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X462 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X463 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X464 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X465 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X466 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X467 a_22404_n7948# VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X468 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X469 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X470 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X471 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X472 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X473 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X474 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X475 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X476 a_13371_n11522# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X477 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X478 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X479 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X480 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X481 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X482 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X483 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X484 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X485 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X486 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X487 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X488 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X489 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X490 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X491 VB2 VB1 a_13371_n10774# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X492 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X493 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X494 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X495 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X496 a_15113_n12143# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X497 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X498 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X499 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X500 a_21723_n12663# IREF IREF AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X501 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X502 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X503 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X504 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X505 dda_0.SUM_N VB3 VO2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X506 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X507 AVSS VB2 a_21723_n13135# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X508 VB1 VB1 a_15113_n13704# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X509 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X510 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X511 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X512 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X513 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X514 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X515 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X516 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X517 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X518 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X519 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X520 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X521 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X522 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X523 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X524 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X525 a_16855_n12608# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X526 dda_0.VD1 VO1 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X527 dda_0.SUM_P VB3 VO1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X528 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X529 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X530 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X531 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X532 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X533 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X534 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X535 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X536 dda_0.VCMFB VCM dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X537 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X538 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X539 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X540 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X541 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
D0 AVSS VO2 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X542 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X543 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X544 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X545 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X546 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X547 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X548 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X549 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X550 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X551 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X552 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X553 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X554 dda_0.VIT_N1 VO1 dda_0.VD1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X555 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X556 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X557 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X558 a_23429_n12663# IREF IREF AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X559 a_13371_n7762# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X560 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X561 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X562 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X563 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X564 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X565 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X566 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X567 AVSS VB2 a_23429_n13135# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X568 a_13887_n10153# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X569 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X570 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X571 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X572 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X573 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X574 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X575 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X576 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X577 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X578 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X579 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X580 a_16339_n11522# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X581 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X582 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X583 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X584 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X585 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X586 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X587 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X588 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X589 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X590 dda_0.VIT_N1 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X591 dda_0.SUM_N VB3 VO2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X592 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X593 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X594 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X595 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X596 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X597 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X598 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X599 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X600 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X601 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X602 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X603 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X604 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X605 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X606 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X607 VB2 VB1 a_15113_n15827# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X608 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X609 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X610 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X611 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X612 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X613 VB2 VB1 a_16339_n15210# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X614 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X615 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X616 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X617 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X618 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X619 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X620 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X621 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X622 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X623 a_15629_n16714# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X624 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X625 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X626 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X627 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X628 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X629 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X630 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X631 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X632 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X633 AVDD VB1 a_13887_n12143# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X634 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X635 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X636 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X637 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X638 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X639 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X640 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X641 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X642 VB1 VB1 a_13371_n13704# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X643 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X644 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X645 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X646 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X647 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X648 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X649 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X650 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X651 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X652 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X653 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X654 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X655 AVDD VB1 a_15629_n12608# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X656 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X657 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X658 AVDD VB1 a_16855_n10774# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X659 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X660 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X661 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X662 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X663 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X664 a_16855_n8649# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X665 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X666 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X667 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X668 a_20870_n12663# VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X669 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X670 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X671 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X672 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X673 a_20017_n12663# IREF IREF AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X674 AVDD VB1 a_14597_n17331# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X675 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X676 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X677 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X678 dda_0.VIT_N2 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X679 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X680 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X681 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X682 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X683 dda_0.SUM_P VB3 VO1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X684 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X685 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X686 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X687 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X688 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X689 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X690 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X691 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X692 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X693 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X694 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X695 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X696 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X697 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X698 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X699 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X700 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X701 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X702 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X703 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X704 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X705 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X706 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X707 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X708 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X709 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X710 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X711 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X712 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X713 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X714 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X715 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X716 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X717 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X718 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X719 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X720 VB3 VB1 a_13371_n15827# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X721 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X722 a_22576_n12663# VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X723 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X724 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X725 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X726 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X727 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X728 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X729 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X730 dda_0.VD2 VO2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X731 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X732 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X733 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X734 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X735 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X736 VO2 VB3 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X737 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X738 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X739 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X740 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X741 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X742 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X743 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X744 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X745 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X746 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X747 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X748 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X749 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X750 a_14597_n10774# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X751 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X752 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X753 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X754 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X755 AVSS VB2 a_20017_n13135# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X756 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X757 a_15113_n11522# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X758 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X759 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X760 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X761 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X762 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X763 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X764 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X765 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X766 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X767 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X768 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X769 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X770 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X771 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X772 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X773 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X774 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X775 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X776 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X777 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X778 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X779 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X780 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X781 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X782 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X783 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X784 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X785 AVDD VB1 a_16855_n7762# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X786 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X787 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X788 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X789 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X790 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X791 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X792 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X793 AVDD VB1 a_13887_n8649# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X794 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X795 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X796 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X797 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X798 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X799 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X800 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X801 AVDD VB1 a_16855_n13704# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X802 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X803 a_15629_n13237# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X804 VB2 VB1 a_15113_n10153# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X805 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X806 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X807 a_13887_n17331# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X808 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X809 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X810 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X811 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X812 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X813 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X814 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X815 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X816 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X817 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X818 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X819 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X820 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X821 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X822 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X823 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X824 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X825 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X826 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X827 AVDD VB1 a_14597_n8649# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X828 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X829 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X830 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X831 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X832 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X833 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X834 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X835 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X836 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X837 dda_0.VIT_N2 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X838 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X839 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X840 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X841 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X842 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X843 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X844 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X845 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X846 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X847 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X848 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X849 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X850 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X851 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X852 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X853 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X854 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X855 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X856 a_13371_n15210# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X857 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X858 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X859 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X860 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X861 a_21723_n13135# VB2 VB2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X862 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X863 VB2 VB1 a_16339_n16714# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X864 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X865 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X866 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X867 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X868 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X869 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X870 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X871 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X872 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X873 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X874 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X875 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X876 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X877 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X878 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X879 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X880 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X881 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X882 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X883 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X884 AVDD VB1 a_16855_n15827# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X885 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X886 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X887 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X888 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X889 AVDD VB1 a_13887_n11522# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X890 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X891 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X892 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X893 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X894 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X895 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X896 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X897 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X898 a_14597_n13704# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X899 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X900 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X901 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X902 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X903 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X904 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X905 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X906 VO1 VB3 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X907 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X908 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X909 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X910 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X911 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X912 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X913 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X914 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X915 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X916 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X917 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X918 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X919 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X920 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X921 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X922 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X923 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X924 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X925 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X926 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X927 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X928 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X929 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X930 a_23429_n13135# VB2 VB2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X931 VB3 VB1 a_13371_n10153# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X932 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X933 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X934 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X935 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X936 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X937 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X938 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X939 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X940 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X941 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X942 a_15113_n7762# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X943 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X944 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X945 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X946 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X947 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X948 dda_0.VIT_N2 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X949 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X950 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X951 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X952 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X953 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X954 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X955 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X956 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X957 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X958 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X959 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X960 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X961 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X962 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X963 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X964 dda_0.VCMFB VCM dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X965 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X966 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X967 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X968 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X969 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X970 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X971 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X972 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X973 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X974 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X975 a_16339_n15210# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X976 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X977 dda_0.SUM_N VB3 VO2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X978 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X979 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X980 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X981 dda_0.VIT_N2 VO2 dda_0.VD2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X982 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X983 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X984 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X985 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X986 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X987 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X988 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X989 a_14597_n15827# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X990 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X991 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X992 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X993 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X994 AVDD VB1 a_14597_n14323# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X995 dda_0.VIT_N1 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X996 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X997 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X998 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X999 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1000 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1001 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1002 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1003 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1004 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1005 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1006 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1007 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1008 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1009 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1010 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1011 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1012 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1013 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1014 a_15629_n12608# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1015 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1016 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1017 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1018 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1019 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1020 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1021 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1022 dda_0.VD1 VO1 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1023 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1024 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1025 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1026 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1027 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1028 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1029 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1030 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1031 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1032 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1033 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1034 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1035 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1036 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1037 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1038 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1039 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1040 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1041 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1042 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1043 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1044 a_20870_n13135# IREF AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1045 VB2 VB1 a_15113_n17331# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1046 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1047 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1048 a_20017_n13135# VB2 VB2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1049 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1050 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1051 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1052 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1053 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1054 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1055 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1056 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1057 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1058 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1059 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1060 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1061 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1062 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1063 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1064 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1065 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1066 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1067 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1068 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1069 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1070 VB1 VB1 a_16339_n13237# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1071 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1072 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1073 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1074 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1075 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1076 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1077 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1078 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1079 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1080 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1081 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1082 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1083 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1084 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1085 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1086 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1087 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1088 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1089 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1090 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1091 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1092 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1093 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1094 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1095 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1096 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1097 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1098 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1099 AVDD VB1 a_16855_n10153# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1100 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1101 a_22576_n13135# IREF AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1102 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1103 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1104 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1105 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1106 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1107 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1108 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1109 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1110 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1111 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1112 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1113 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1114 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1115 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1116 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1117 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1118 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1119 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1120 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1121 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1122 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1123 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1124 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1125 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1126 dda_0.SUM_N VB3 VO2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1127 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1128 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1129 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1130 dda_0.VD2 VO2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1131 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1132 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1133 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1134 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1135 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1136 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1137 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1138 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1139 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1140 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1141 a_13887_n14323# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1142 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1143 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1144 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1145 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1146 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1147 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1148 a_13371_n16714# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1149 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1150 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1151 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1152 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1153 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1154 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1155 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1156 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1157 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1158 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1159 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1160 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1161 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1162 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1163 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1164 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1165 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1166 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1167 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1168 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1169 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1170 a_15113_n15210# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1171 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1172 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1173 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1174 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1175 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1176 VB3 VB1 a_13371_n17331# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1177 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1178 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1179 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1180 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1181 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1182 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1183 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1184 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1185 dda_0.SUM_P VB3 VO1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1186 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1187 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1188 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1189 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1190 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1191 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1192 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1193 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1194 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1195 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1196 a_14597_n10153# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1197 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1198 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1199 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1200 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1201 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1202 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1203 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1204 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1205 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1206 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1207 VB4 VB4 a_22662_n7484# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1208 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1209 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1210 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1211 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1212 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1213 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1214 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1215 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1216 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1217 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1218 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1219 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1220 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1221 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1222 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1223 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1224 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1225 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1226 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1227 VB1 IREF a_20870_n14041# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1228 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1229 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1230 dda_0.VCMFB VCM dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1231 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1232 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1233 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1234 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1235 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1236 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1237 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1238 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1239 a_16339_n16714# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1240 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1241 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1242 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1243 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1244 dda_0.VIT_N1 VO1 dda_0.VD1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1245 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1246 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1247 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1248 AVDD VB1 a_14597_n12143# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1249 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1250 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1251 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1252 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1253 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1254 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1255 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1256 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1257 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1258 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1259 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1260 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1261 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1262 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1263 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1264 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1265 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1266 VB4 VB2 a_20870_n11758# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1267 VB1 VB1 a_16339_n12608# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1268 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1269 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1270 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1271 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1272 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1273 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1274 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1275 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1276 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1277 AVDD VB1 a_13887_n15210# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1278 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1279 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1280 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1281 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1282 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1283 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1284 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1285 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1286 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1287 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1288 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1289 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1290 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1291 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1292 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1293 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1294 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1295 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1296 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1297 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1298 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1299 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1300 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1301 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1302 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1303 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1304 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1305 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1306 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1307 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1308 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1309 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1310 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1311 VB2 VB1 a_15113_n8649# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1312 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1313 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1314 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1315 a_13371_n13237# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1316 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1317 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1318 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1319 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1320 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1321 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1322 AVDD VB1 a_16855_n17331# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1323 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1324 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1325 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1326 dda_0.SUM_P VB3 VO1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1327 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1328 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1329 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1330 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1331 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1332 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1333 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1334 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1335 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1336 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1337 VO2 VB3 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1338 VB4 VB4 a_22662_n7948# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1339 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1340 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1341 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1342 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1343 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1344 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1345 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1346 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1347 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1348 VB2 VB1 a_15113_n14323# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1349 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1350 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1351 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1352 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1353 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1354 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1355 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1356 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1357 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1358 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1359 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1360 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1361 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1362 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1363 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1364 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1365 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1366 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1367 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1368 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1369 a_13887_n12143# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1370 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1371 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1372 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1373 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1374 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1375 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1376 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1377 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1378 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1379 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1380 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1381 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1382 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1383 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1384 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1385 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1386 dda_0.VD2 VO2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1387 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1388 VO1 VB3 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1389 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1390 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1391 a_16855_n10774# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1392 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1393 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1394 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1395 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1396 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1397 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1398 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1399 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1400 a_15113_n16714# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1401 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1402 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1403 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1404 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1405 a_14597_n17331# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1406 a_16339_n13237# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1407 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1408 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1409 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1410 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1411 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1412 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1413 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1414 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1415 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1416 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1417 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1418 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1419 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1420 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1421 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1422 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1423 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1424 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1425 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1426 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1427 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1428 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1429 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1430 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1431 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1432 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1433 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1434 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1435 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1436 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1437 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1438 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1439 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1440 a_23540_n15948# VB3 a_23282_n15948# AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1441 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1442 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1443 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1444 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1445 a_13371_n8649# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1446 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1447 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1448 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1449 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1450 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1451 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1452 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1453 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1454 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1455 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1456 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1457 VB3 VB1 a_13371_n14323# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1458 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1459 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1460 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1461 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1462 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1463 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1464 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1465 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1466 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1467 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1468 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1469 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1470 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1471 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1472 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1473 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1474 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1475 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1476 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1477 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1478 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1479 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1480 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1481 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1482 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1483 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1484 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1485 AVDD VB1 a_14597_n11522# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1486 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1487 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1488 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1489 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1490 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1491 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1492 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1493 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1494 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1495 a_13371_n12608# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1496 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1497 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1498 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1499 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1500 AVDD VB1 a_15629_n10774# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1501 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1502 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1503 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1504 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1505 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1506 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1507 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1508 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1509 AVDD VB1 a_13887_n16714# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1510 a_16855_n13704# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1511 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1512 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1513 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1514 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1515 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1516 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1517 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1518 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1519 dda_0.VIT_N2 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1520 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1521 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1522 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1523 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1524 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1525 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1526 AVDD VB1 a_15629_n9266# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1527 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1528 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1529 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1530 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1531 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1532 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1533 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1534 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1535 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1536 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1537 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1538 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1539 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1540 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1541 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1542 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1543 VB2 VB1 a_16339_n9266# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1544 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1545 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1546 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1547 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1548 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1549 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1550 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1551 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1552 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1553 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1554 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1555 a_15113_n13237# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1556 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1557 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1558 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1559 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1560 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1561 VB1 VB1 a_15113_n12143# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1562 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1563 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1564 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1565 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1566 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1567 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1568 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1569 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1570 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1571 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1572 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1573 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1574 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1575 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1576 a_16339_n12608# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1577 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1578 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1579 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1580 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1581 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1582 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1583 a_16855_n15827# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1584 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1585 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1586 a_13887_n11522# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1587 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1588 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1589 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1590 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1591 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1592 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1593 AVDD VB1 a_16855_n14323# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1594 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1595 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1596 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1597 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1598 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1599 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1600 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1601 dda_0.VIT_N1 VO1 dda_0.VD1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1602 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1603 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1604 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1605 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1606 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1607 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1608 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1609 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1610 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1611 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1612 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1613 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1614 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1615 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1616 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1617 AVDD VB1 a_15629_n13704# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1618 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1619 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1620 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1621 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1622 dda_0.VIT_N1 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1623 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1624 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1625 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1626 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1627 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1628 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1629 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1630 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1631 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1632 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1633 AVDD VB1 a_16855_n8649# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1634 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1635 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1636 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1637 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1638 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1639 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1640 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1641 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1642 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1643 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1644 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1645 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1646 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1647 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1648 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1649 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1650 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1651 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1652 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1653 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1654 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1655 a_15629_n9266# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1656 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1657 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1658 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1659 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1660 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1661 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1662 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1663 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1664 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1665 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1666 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1667 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1668 a_13887_n9266# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1669 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1670 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1671 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1672 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1673 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1674 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1675 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1676 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1677 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1678 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1679 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1680 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1681 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1682 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1683 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1684 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1685 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1686 a_16339_n9266# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1687 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1688 AVDD VB1 a_13887_n13237# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1689 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1690 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1691 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1692 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1693 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1694 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1695 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1696 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1697 VB1 VB1 a_13371_n12143# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1698 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1699 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1700 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1701 a_14597_n14323# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1702 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1703 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1704 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1705 a_14597_n9266# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1706 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1707 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1708 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1709 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1710 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
D1 AVSS VI_1A sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X1711 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1712 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1713 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1714 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
D2 AVSS VI_2B sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X1715 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1716 dda_0.VIT_N2 VO2 dda_0.VD2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1717 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1718 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1719 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1720 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1721 AVDD VB1 a_15629_n15827# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1722 dda_0.SUM_N VB3 VO2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1723 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1724 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1725 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1726 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1727 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1728 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1729 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1730 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1731 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1732 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1733 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1734 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1735 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1736 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1737 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1738 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1739 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1740 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1741 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1742 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1743 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1744 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1745 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1746 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1747 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1748 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1749 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1750 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1751 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1752 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1753 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1754 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1755 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1756 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1757 a_15113_n12608# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1758 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1759 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1760 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1761 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1762 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1763 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1764 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1765 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1766 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1767 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1768 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1769 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1770 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1771 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1772 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1773 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1774 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1775 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1776 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1777 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1778 a_16855_n10153# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1779 a_22662_n8251# VB4 a_22404_n8251# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1780 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1781 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1782 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1783 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1784 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1785 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1786 a_15113_n8649# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1787 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1788 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1789 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1790 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1791 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1792 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1793 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1794 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1795 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1796 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1797 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1798 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
D3 AVSS VI_1B sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X1799 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1800 VB2 VB1 a_13371_n9266# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1801 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1802 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
D4 AVSS VI_2A sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X1803 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1804 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1805 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1806 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1807 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1808 VB1 VB1 a_15113_n11522# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1809 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1810 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1811 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1812 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1813 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1814 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1815 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1816 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1817 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1818 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1819 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1820 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1821 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1822 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1823 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1824 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1825 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1826 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1827 dda_0.VIT_N1 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1828 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1829 a_15629_n10774# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1830 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1831 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1832 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1833 AVDD VB1 a_14597_n15210# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1834 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1835 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1836 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1837 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1838 AVDD VB1 a_16855_n12143# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1839 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1840 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1841 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1842 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1843 dda_0.VD2 VO2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1844 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1845 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1846 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1847 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1848 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1849 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1850 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1851 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1852 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1853 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1854 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1855 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1856 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1857 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1858 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1859 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1860 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1861 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1862 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1863 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1864 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1865 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1866 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1867 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1868 dda_0.SUM_P VB3 VO1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1869 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1870 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1871 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1872 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1873 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1874 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1875 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1876 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1877 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1878 AVDD VB1 a_13887_n12608# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1879 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1880 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1881 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1882 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1883 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1884 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1885 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1886 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1887 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1888 dda_0.VD1 VO1 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1889 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1890 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1891 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1892 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1893 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1894 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1895 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1896 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1897 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1898 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1899 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1900 AVDD VB1 a_15629_n10153# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1901 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1902 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1903 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1904 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1905 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1906 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1907 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1908 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1909 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1910 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1911 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1912 a_22404_n8251# VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1913 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1914 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1915 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1916 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1917 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1918 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1919 a_22662_n8715# VB4 a_22404_n8715# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1920 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1921 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1922 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1923 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1924 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1925 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1926 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1927 dda_0.VCMFB VCM dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1928 VO2 VB3 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1929 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1930 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1931 dda_0.VD2 VO2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1932 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1933 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1934 a_14597_n12143# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1935 VB1 VB1 a_13371_n11522# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1936 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1937 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1938 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1939 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1940 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1941 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1942 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1943 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1944 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1945 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1946 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1947 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1948 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1949 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1950 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1951 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1952 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1953 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1954 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1955 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1956 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1957 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1958 a_13887_n15210# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1959 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1960 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1961 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1962 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1963 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1964 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1965 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1966 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1967 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1968 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1969 a_15629_n13704# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1970 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1971 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1972 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1973 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1974 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1975 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1976 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1977 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1978 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1979 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1980 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1981 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1982 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1983 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1984 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1985 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1986 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1987 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1988 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1989 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1990 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1991 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1992 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1993 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1994 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1995 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1996 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1997 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X1998 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X1999 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2000 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2001 a_16855_n17331# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2002 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2003 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2004 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2005 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2006 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2007 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2008 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2009 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2010 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2011 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2012 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2013 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2014 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2015 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2016 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2017 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2018 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2019 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2020 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2021 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2022 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2023 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2024 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2025 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2026 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2027 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2028 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2029 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2030 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2031 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2032 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2033 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2034 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2035 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2036 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2037 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2038 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2039 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2040 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2041 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2042 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2043 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2044 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2045 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2046 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2047 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2048 a_15629_n15827# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2049 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2050 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2051 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2052 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2053 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2054 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2055 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2056 a_22404_n8715# VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2057 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2058 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2059 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2060 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2061 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2062 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2063 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2064 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2065 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2066 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2067 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2068 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2069 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2070 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2071 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2072 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2073 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2074 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2075 AVDD VB1 a_15629_n7762# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2076 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2077 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2078 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2079 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2080 VB2 VB1 a_16339_n10774# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2081 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2082 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2083 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2084 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2085 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2086 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2087 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2088 AVDD VB1 a_16855_n11522# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2089 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2090 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2091 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2092 AVDD VB1 a_14597_n16714# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2093 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2094 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2095 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2096 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2097 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2098 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2099 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2100 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2101 VB2 VB1 a_16339_n7762# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2102 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2103 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2104 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2105 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2106 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2107 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2108 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2109 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2110 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2111 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2112 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2113 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2114 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2115 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2116 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2117 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2118 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2119 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2120 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2121 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2122 VB2 VB2 a_20870_n12663# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2123 dda_0.VIT_N2 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2124 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2125 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2126 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2127 AVDD VB1 a_15629_n17331# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2128 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2129 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2130 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2131 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2132 a_23282_n15948# VB3 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2133 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2134 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2135 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2136 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2137 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2138 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2139 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2140 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2141 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2142 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2143 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2144 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2145 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2146 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2147 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2148 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2149 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2150 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2151 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2152 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2153 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2154 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2155 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2156 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2157 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2158 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2159 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2160 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2161 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2162 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2163 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2164 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2165 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2166 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2167 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2168 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2169 a_14597_n11522# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2170 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2171 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2172 VB3 VB1 a_15113_n15210# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2173 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2174 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2175 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2176 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2177 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2178 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2179 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2180 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2181 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2182 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2183 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2184 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2185 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2186 dda_0.SUM_N VB3 VO2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2187 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2188 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2189 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2190 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2191 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2192 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
D5 AVSS IREF sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X2193 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2194 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2195 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2196 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2197 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2198 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2199 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2200 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2201 a_15629_n7762# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2202 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2203 a_13887_n16714# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2204 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2205 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2206 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2207 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2208 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2209 VB1 VB1 a_16339_n13704# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2210 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2211 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2212 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2213 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2214 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2215 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2216 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2217 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2218 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2219 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2220 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2221 a_13887_n7762# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2222 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2223 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2224 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2225 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2226 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2227 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2228 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2229 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2230 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2231 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2232 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2233 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2234 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2235 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2236 a_16339_n7762# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2237 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2238 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2239 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2240 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2241 a_15629_n10153# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2242 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2243 a_14597_n7762# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2244 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2245 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2246 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2247 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2248 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2249 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2250 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2251 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2252 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2253 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2254 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2255 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2256 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2257 VO1 VB3 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2258 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2259 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2260 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2261 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2262 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2263 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2264 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2265 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2266 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2267 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2268 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2269 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2270 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2271 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2272 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2273 AVDD VB1 a_14597_n13237# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2274 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2275 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2276 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2277 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2278 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2279 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2280 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2281 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2282 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2283 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2284 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2285 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2286 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2287 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2288 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2289 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2290 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2291 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2292 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2293 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2294 dda_0.SUM_N VB3 VO2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2295 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2296 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2297 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2298 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2299 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2300 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2301 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2302 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2303 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2304 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2305 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2306 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2307 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2308 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2309 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2310 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2311 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2312 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2313 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2314 VB3 VB1 a_16339_n15827# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
D6 AVSS VO1 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X2315 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2316 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2317 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2318 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2319 VB2 VB1 a_13371_n15210# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2320 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2321 a_16855_n14323# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2322 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2323 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2324 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2325 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2326 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2327 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2328 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2329 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2330 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2331 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2332 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2333 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2334 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2335 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2336 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2337 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2338 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2339 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2340 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2341 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2342 a_13371_n10774# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2343 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2344 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2345 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2346 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2347 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2348 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2349 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2350 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2351 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2352 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2353 dda_0.VIT_N2 VO2 dda_0.VD2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2354 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2355 dda_0.SUM_P VB3 VO1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2356 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2357 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2358 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2359 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2360 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2361 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2362 VB1 IREF a_22576_n14041# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2363 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2364 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2365 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2366 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2367 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2368 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2369 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2370 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2371 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2372 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2373 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2374 VB2 VB1 a_13371_n7762# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2375 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2376 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2377 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2378 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2379 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2380 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2381 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2382 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2383 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2384 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2385 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2386 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2387 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2388 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2389 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2390 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2391 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2392 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2393 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2394 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2395 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2396 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2397 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2398 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2399 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2400 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2401 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2402 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2403 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2404 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2405 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2406 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2407 a_22662_n9018# VB4 a_22404_n9018# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2408 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2409 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2410 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2411 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2412 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2413 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2414 a_13887_n13237# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2415 dda_0.VIT_N1 VO1 dda_0.VD1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2416 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2417 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2418 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2419 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2420 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2421 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2422 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2423 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2424 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2425 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2426 dda_0.VCMFB VCM dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2427 VB4 VB2 a_22576_n11758# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2428 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2429 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2430 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2431 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2432 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2433 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2434 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2435 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2436 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2437 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2438 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2439 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2440 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2441 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2442 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2443 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2444 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2445 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2446 a_16339_n10774# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2447 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2448 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2449 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2450 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2451 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2452 AVDD VB1 a_15629_n14323# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2453 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2454 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2455 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2456 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2457 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2458 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2459 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2460 VB3 VB1 a_15113_n16714# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2461 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2462 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2463 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2464 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2465 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2466 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2467 dda_0.VCMFB VCM dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2468 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2469 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2470 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2471 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2472 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2473 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2474 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2475 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2476 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2477 AVDD VB1 a_16855_n15210# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2478 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2479 a_13371_n13704# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2480 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2481 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2482 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2483 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2484 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2485 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2486 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2487 dda_0.VD1 VO1 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2488 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2489 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2490 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2491 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2492 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2493 IREF IREF a_20870_n13135# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2494 a_15629_n17331# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2495 AVDD VB1 a_14597_n12608# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2496 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2497 dda_0.VIT_N2 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2498 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2499 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2500 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2501 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2502 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2503 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2504 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2505 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2506 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2507 VB3 VB1 a_16339_n10153# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2508 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2509 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2510 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2511 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2512 dda_0.VIT_N1 VO1 dda_0.VD1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2513 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2514 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2515 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2516 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2517 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2518 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2519 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2520 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2521 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2522 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2523 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2524 AVSS VB2 a_21723_n14041# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2525 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2526 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2527 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2528 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2529 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2530 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2531 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2532 a_16855_n9266# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2533 dda_0.VCMFB VCM dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2534 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2535 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2536 a_22404_n9018# VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2537 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2538 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2539 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2540 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2541 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2542 VB3 VB3 a_23798_n15948# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2543 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2544 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2545 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2546 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2547 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2548 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2549 a_13371_n15827# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2550 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2551 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2552 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2553 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2554 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2555 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2556 a_14597_n15210# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2557 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2558 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2559 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2560 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2561 a_16855_n12143# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2562 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2563 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2564 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2565 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2566 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2567 VB2 VB1 a_13371_n16714# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2568 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2569 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2570 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2571 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2572 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2573 a_16339_n13704# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2574 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2575 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2576 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2577 AVSS VB2 a_23429_n14041# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2578 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2579 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2580 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2581 AVSS IREF a_21723_n11758# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2582 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2583 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2584 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2585 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2586 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2587 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2588 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2589 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2590 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2591 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2592 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2593 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2594 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2595 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2596 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2597 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2598 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2599 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2600 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2601 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2602 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2603 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2604 a_13887_n12608# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2605 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2606 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2607 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2608 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2609 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2610 a_15113_n10774# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2611 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2612 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2613 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2614 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2615 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2616 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2617 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2618 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2619 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2620 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2621 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2622 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2623 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2624 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2625 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2626 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2627 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2628 dda_0.VCMFB VCM dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2629 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2630 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2631 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2632 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2633 AVSS IREF a_23429_n11758# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2634 VB1 VB1 a_15113_n13237# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2635 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2636 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2637 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2638 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2639 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2640 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2641 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2642 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2643 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2644 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2645 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2646 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2647 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2648 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2649 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2650 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2651 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2652 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2653 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2654 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2655 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2656 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2657 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2658 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2659 AVDD VB1 a_13887_n9266# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2660 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2661 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2662 a_16339_n15827# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2663 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2664 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2665 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2666 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2667 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2668 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2669 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2670 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2671 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2672 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2673 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2674 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2675 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2676 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2677 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2678 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2679 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2680 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2681 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2682 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2683 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2684 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2685 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2686 AVDD VB1 a_14597_n9266# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2687 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2688 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2689 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2690 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2691 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2692 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2693 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2694 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2695 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2696 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2697 AVDD VB1 a_15629_n12143# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2698 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2699 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2700 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2701 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2702 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2703 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2704 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2705 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2706 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2707 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2708 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2709 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2710 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2711 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2712 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2713 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2714 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2715 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2716 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2717 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2718 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2719 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2720 AVSS VB2 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2721 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2722 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2723 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2724 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2725 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2726 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2727 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2728 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2729 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2730 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2731 dda_0.VD2 VO2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2732 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2733 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2734 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2735 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2736 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2737 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2738 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2739 AVDD VB1 a_16855_n16714# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2740 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2741 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2742 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2743 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2744 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2745 VB3 VB1 a_16339_n17331# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2746 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2747 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2748 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2749 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2750 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2751 AVDD VB1 a_13887_n10774# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2752 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2753 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2754 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2755 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2756 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2757 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2758 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2759 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2760 a_15113_n13704# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2761 VB1 VB1 a_13371_n13237# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2762 a_13371_n10153# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2763 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2764 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2765 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2766 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2767 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2768 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2769 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2770 AVSS VB2 a_20017_n14041# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2771 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2772 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2773 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2774 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2775 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2776 VB4 VB4 a_22662_n8251# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2777 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2778 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2779 dda_0.SUM_P VB3 VO1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2780 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2781 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2782 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2783 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2784 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2785 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2786 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2787 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2788 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2789 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2790 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2791 a_15629_n14323# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2792 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2793 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2794 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2795 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2796 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2797 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2798 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2799 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2800 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2801 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2802 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2803 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2804 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2805 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2806 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2807 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2808 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2809 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2810 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2811 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2812 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2813 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2814 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2815 AVSS IREF a_20017_n11758# AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2816 a_16855_n11522# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2817 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2818 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2819 a_14597_n16714# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2820 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2821 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2822 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2823 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2824 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2825 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2826 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2827 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2828 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2829 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2830 VO2 VB3 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2831 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2832 a_15113_n15827# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2833 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2834 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2835 VB1 VB1 a_15113_n12608# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2836 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2837 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2838 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2839 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2840 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2841 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2842 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2843 VO1 VB3 dda_0.SUM_P AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2844 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2845 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2846 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2847 a_16339_n10153# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2848 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2849 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2850 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2851 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2852 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2853 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2854 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2855 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2856 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2857 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2858 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2859 a_21723_n14041# VB2 VB4 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2860 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2861 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2862 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2863 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2864 AVDD VB1 a_13887_n13704# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2865 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2866 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2867 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2868 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2869 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2870 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2871 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2872 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2873 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2874 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2875 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2876 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2877 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2878 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2879 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2880 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2881 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2882 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2883 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2884 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2885 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2886 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2887 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2888 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2889 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2890 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2891 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2892 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2893 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2894 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2895 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2896 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2897 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2898 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2899 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2900 VO2 VB3 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2901 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2902 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2903 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2904 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2905 AVSS VB2 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2906 AVDD VB1 a_16855_n13237# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2907 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2908 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2909 VB4 VB4 a_22662_n8715# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2910 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2911 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2912 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2913 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2914 dda_0.VIT_N2 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2915 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2916 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2917 a_23429_n14041# VB2 VB4 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2918 a_21723_n11758# IREF VB1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2919 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2920 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2921 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2922 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2923 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2924 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2925 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2926 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2927 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2928 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2929 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2930 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2931 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2932 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2933 AVDD VB1 a_15629_n11522# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2934 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2935 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2936 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2937 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2938 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2939 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2940 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2941 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2942 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2943 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2944 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2945 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2946 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2947 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2948 VB1 VB1 a_13371_n12608# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2949 AVDD VB1 a_13887_n15827# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2950 AVDD VB1 a_15629_n8649# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2951 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2952 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2953 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2954 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2955 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2956 AVDD dda_0.VD2 dda_0.VD2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2957 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2958 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2959 dda_0.VIT_N1 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2960 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2961 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2962 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2963 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2964 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2965 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2966 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2967 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2968 a_13371_n17331# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2969 a_23429_n11758# IREF VB1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2970 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2971 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2972 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2973 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2974 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2975 VB3 VB1 a_16339_n8649# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2976 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2977 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2978 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2979 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2980 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2981 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2982 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2983 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2984 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2985 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2986 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2987 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2988 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2989 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2990 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2991 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2992 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2993 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2994 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2995 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2996 a_14597_n13237# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2997 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2998 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2999 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3000 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3001 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3002 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3003 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3004 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3005 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3006 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3007 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3008 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3009 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3010 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3011 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3012 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3013 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3014 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3015 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3016 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3017 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3018 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3019 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3020 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3021 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3022 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3023 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3024 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3025 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3026 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3027 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3028 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3029 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3030 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3031 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3032 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3033 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3034 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3035 a_20870_n14041# IREF AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3036 a_15113_n10153# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3037 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3038 a_20017_n14041# VB2 VB4 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3039 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3040 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3041 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3042 a_15629_n12143# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3043 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3044 VB3 VB1 a_16339_n14323# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3045 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3046 dda_0.VCMFB VCM dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3047 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3048 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3049 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3050 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3051 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3052 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3053 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3054 dda_0.VIT_N2 VO2 dda_0.VD2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3055 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3056 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3057 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3058 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3059 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3060 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3061 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3062 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3063 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3064 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3065 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3066 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3067 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3068 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3069 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3070 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3071 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3072 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3073 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3074 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3075 dda_0.VIT_N1 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3076 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3077 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3078 AVSS VB2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3079 a_16339_n17331# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3080 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3081 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3082 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3083 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3084 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3085 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3086 a_22576_n14041# IREF AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3087 a_20870_n11758# VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3088 a_20017_n11758# IREF VB1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3089 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3090 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3091 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3092 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3093 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3094 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3095 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3096 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3097 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
D7 AVSS VCM sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X3098 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3099 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3100 a_15629_n8649# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3101 a_16855_n7762# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3102 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3103 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3104 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3105 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3106 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3107 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3108 dda_0.VD1 VO1 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3109 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3110 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3111 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3112 a_13887_n8649# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3113 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3114 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3115 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3116 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3117 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3118 AVDD VB1 a_16855_n12608# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3119 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3120 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3121 AVDD dda_0.VCMFB dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3122 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3123 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3124 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3125 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3126 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3127 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3128 AVSS VB2 dda_0.SUM_N AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3129 a_16339_n8649# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3130 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3131 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3132 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3133 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3134 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3135 a_14597_n8649# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3136 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3137 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3138 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3139 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3140 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3141 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3142 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3143 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3144 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3145 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3146 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3147 a_22576_n11758# VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3148 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3149 dda_0.VCMFB VCM dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3150 dda_0.VIT_N1 VCM dda_0.VCMFB AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3151 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3152 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3153 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3154 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3155 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3156 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3157 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3158 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3159 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3160 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3161 AVDD VB1 a_13887_n10153# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3162 VB3 VB1 a_15113_n9266# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3163 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3164 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3165 dda_0.SUM_P VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3166 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3167 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3168 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3169 dda_0.SUM_P VI_2B dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3170 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3171 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3172 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3173 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3174 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3175 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3176 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3177 dda_0.VIT_N1 VO1 dda_0.VD1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3178 dda_0.VD6 VB4 VO2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3179 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3180 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3181 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3182 VO1 VB4 dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3183 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3184 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3185 dda_0.VD2 dda_0.VD2 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3186 dda_0.VD6 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3187 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3188 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3189 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3190 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3191 dda_0.VD2 VO2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3192 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3193 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3194 a_16855_n15210# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3195 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3196 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3197 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3198 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3199 dda_0.VCMFB VCM dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3200 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3201 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3202 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3203 dda_0.SUM_P VI_1A dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3204 dda_0.SUM_N VI_1B dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3205 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3206 dda_0.VIT_N2 VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3207 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3208 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3209 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3210 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3211 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3212 a_14597_n12608# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3213 dda_0.VD2 VO2 dda_0.VIT_N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3214 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3215 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3216 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3217 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3218 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3219 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3220 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3221 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3222 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3223 dda_0.VD1 dda_0.VD1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3224 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3225 AVDD VB1 a_13887_n7762# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3226 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3227 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3228 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3229 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3230 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3231 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3232 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3233 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3234 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3235 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3236 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3237 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3238 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3239 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3240 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3241 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3242 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3243 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3244 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3245 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3246 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3247 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3248 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3249 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3250 VB3 VB1 a_13371_n8649# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3251 AVDD VB1 a_14597_n7762# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3252 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3253 AVDD dda_0.VD1 dda_0.VD1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3254 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3255 dda_0.VD5 VB4 VO1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3256 VO2 VB4 dda_0.VD6 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3257 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3258 dda_0.VD1 VO1 dda_0.VIT_N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3259 dda_0.SUM_P VB3 VO1 AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3260 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3261 a_15113_n17331# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3262 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3263 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3264 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3265 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3266 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3267 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3268 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3269 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3270 dda_0.VIT_P2 VI_2A dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3271 a_23798_n15948# VB3 a_23540_n15948# AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3272 AVDD VB1 dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3273 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3274 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3275 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3276 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3277 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3278 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3279 dda_0.VIT_P1 VI_1B dda_0.SUM_N AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3280 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3281 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3282 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3283 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3284 dda_0.SUM_N VB2 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3285 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3286 dda_0.VD5 dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3287 dda_0.VIT_P1 VI_1A dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3288 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3289 dda_0.VIT_P2 VI_2B dda_0.SUM_P AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3290 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3291 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3292 a_13371_n14323# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3293 dda_0.VIT_P1 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3294 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3295 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3296 VB1 VB1 a_16339_n12143# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3297 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3298 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3299 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3300 a_15629_n11522# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3301 dda_0.SUM_N VI_2A dda_0.VIT_P2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3302 dda_0.VCMFB dda_0.VCMFB AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3303 AVDD dda_0.VCMFB dda_0.VCMFB AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3304 AVDD dda_0.VCMFB dda_0.VD5 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3305 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3306 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3307 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3308 AVDD VB1 dda_0.VIT_P1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3309 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3310 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3311 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3312 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3313 dda_0.VIT_P2 VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X3314 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3315 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3316 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
.ends

